TEST CIRCUIT
*
*Q1 N001 N002 N003 PNP
*V1 N002 0 SIN(-5 1 10)
*R1 N001 N004 9.5k
*V2 N004 0 -20
*R2 N003 0 3k
*
Q1 N002 N003 N004 PNP
R1 N001 N002 10k
R2 N004 0 3k
V1 N003 0 SINE(-5 1 10)
V2 N001 0 -20
*
.model PNP PNP
.tran 0.0001 0.5 0
.end