TEST CIRCUIT
*
V1 N003 0 SINE(0 5 10)
R1 N004 0 2k
R2 N001 N002 2k
V2 N001 0 -10
M1 N002 N003 N004 0 PMOS
*
.model PNP PNP
.model NPN NPN
.model PMOS PMOS
.model NMOS NMOS
.tran 0.0001 0.5 0
.end
