TEST CIRCUIT
*
* DIFFERENTIAL AMPLIFIER
Q1 N003 N001 N002 0 NPN
Q2 N004 N001 N002 0 PNP
V1 N001 0 SIN(0 1 5)
V2 N004 0 -20
V3 N003 0 20
R1 N002 0 10k
*
.options Gmin=2
*
.model D D
.model PNP PNP
.model NPN NPN
.model NMOS NMOS
.model PMOS PMOS
.tran 0.00001 1 0
.options Gmin=1m
.end
