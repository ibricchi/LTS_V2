Dependent source test
*
V1 N001 0 5
R1 N002 N001 1k
C1 N002 0 1n
R2 N002 0 1k
*
.tran 0.0001 .2 0 1
.end