Dependent source test
*
XU1 N001 N003 N002 Ideal
R1 N002 N001 2k
R2 N001 0 1k
V1 N003 0 20
*
.tran 0.0001 .5 0 1
.end