TEST CIRCUIT
*
M1 N003 N002 0 0 NMOS
M2 N002 N002 0 0 NMOS
I1 0 N002 100m
R1 N001 N003 100
V1 N001 0 36
*
.model PNP PNP
.model NPN NPN
.model NMOS NMOS
.model PMOS PMOS
.tran 0.00001 1 0
.end
