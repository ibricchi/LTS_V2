Simple Diode
*
V1 N1 0 SIN(0 1 10)
R1 N2 0 1k
D1 N1 N2
*
.tran 0.1 1 0 0.00001
.end
