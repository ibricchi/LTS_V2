Inverting Op-Amp from EE1 Term 2 Labs
QT2[3] N012 0 N014 0 2N2907
QT1[3] N016 N001 N014 0 2N2907
QT2[1] N006 N006 N003 0 2N2907
QT1[1] N008 N006 N003 0 2N2907
QT2[2] N014 N008 N006 0 2N2907
R1 N008 N017 8.3k
QT2[4] N012 N016 N017 0 2N2222
QT1[4] N016 N016 N017 0 2N2222
QT2[6] N011 N015 N017 0 2N2222
V-Vcc N017 0 0
QT1[5] N005 N005 N003 0 2N2907
QT2[5] N004 N005 N003 0 2N2907
R2 N005 N017 9.3k
R3 N015 N017 1.5k
QT1[6] N011 N012 N015 0 2N2222
QT1[7] N004 N004 N010 0 2N2222
QT2[7] N003 N004 N007 0 2N2222
QT2[8] N004 N007 N002 0 2N2222
RCL1 N002 N007 2
RCL2 N009 N002 2
QT1[2] N011 N009 N002 0 2N2907
QT1[9] N011 N011 N010 0 2N2907
QT2[9] N017 N011 N009 0 2N2907
V+Vcc N003 0 0
C N011 N012 10p
Vin N013 0 SIN(0 5m 1)
Rf N002 N001 25k
Rin N001 N013 5k
.model 2N2222 NPN (VAF=100 BF=200 BR=3)
.model 2N2907 PNP (VAF=120 BF=250 BR=3)
.tran 10u .5
.options gmin=1p abstol=0.01 imax=1000
.END
