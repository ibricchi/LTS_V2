Simple Diode
*
V1 N1 0 SIN(0 1 10)
R1 N2 0 1
R2 N1 N2 1
*
.tran 0.1 1 0 0.001
.end
