TEST CIRCUIT
*
* DIFFERENTIAL AMPLIFIER
*Q1 N003 N001 N002 0 NPN
*Q2 N004 N001 N002 0 PNP
*V1 N001 0 SIN(0 1 5)
*V2 N004 0 -20
*V3 N003 0 20
*R1 N002 0 10k
*
V1 N001 0 PULSE(2 5 0.1 0.2 0 0.1 0.3)
R2 N001 N003 1k
R1 N003 0 1k
R3 N002 0 2k
F1 N003 N002 V1 2
.tran 10u 1 0
.options Gmin=1p
.end
