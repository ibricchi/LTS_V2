TEST CIRCUIT
*
V1 N001 0 SINE(0 5m 10)
R1 N002 N001 10k
R2 N003 N002 10k
D1 N003 N006
D2 N006 N002
XU1 N002 0 N006
XU2 N004 0 N005 ideal
R3 N003 N004 10k
R4 N005 N004 10k
*
*Q1 N001 N003 N004 0 NPN
*R1 N002 N001 4.7k
*R2 N004 0 1k
*C1 N004 0 20µ
*R3 N003 0 1k
*R4 N002 N003 4.7k
*V2 N002 0 9
*V1 N003 0 Sin(0 2 10)
*
.model PNP PNP
.model NPN NPN
.model NMOS NMOS
.model PMOS PMOS
.tran 0.00001 1 0
.end
